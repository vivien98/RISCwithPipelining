library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity hazard is
	port(clk,shift,wr: in std_logic ;writeData : in std_logic_vector(7 downto 0);bit1: out std_logic);
end entity;
architecture kahipan of hazard is

begin

end kahipan;

